//run_sv2v

`include "ibex_pkg.sv"
import ibex_pkg::*;

module ibex_compressed_decoder_stimulus (
  output  logic        clk_i,
  output  logic        rst_ni,
  output  logic        valid_i,
  output  logic [31:0] instr_i,
  output  logic [15:0] enum_dpi,
);
 
endmodule